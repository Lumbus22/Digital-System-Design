module sp1(x1, x2, x3, F);

input x1, x2, x3;

output F;

assign F = (~x2 & x3) | (x1 & ~x2) | (~x1 & x2 & x3) | (x1 & ~x3);

endmodule